module rom (
  input wire [6:0] address,
  input wire clk,
  output reg [15:0] data
);


  // Define your ROM contents here
  reg [15:0] rom_contents [0:2**6-1] = {
    // Fill in your data values here
    // 16-bit ROM with 64 address locations
    16'b0000000000011100; 
    16'b0000000000011010;    
    16'b0000000000010100;    
    16'b0000000000000110;    
    16'b1111111111110001;    
    16'b1111111111010110;    
    16'b1111111110111011;    
    16'b1111111110100111;    
    16'b1111111110100111;    
    16'b1111111111000011;    
    16'b0000000000000000;    
    16'b0000000001011000;    
    16'b0000000010111010;    
    16'b0000000100001101;    
    16'b0000000100110001;    
    16'b0000000100001001;    
    16'b0000000010000111;    
    16'b1111111110110000;    
    16'b1111111010100100;    
    16'b1111110110011010;    
    16'b1111110011011110;    
    16'b1111110010111100;    
    16'b1111110101110111;    
    16'b1111111100110011;    
    16'b0000000111101010;    
    16'b0000010101100111;    
    16'b0000100101001011;    
    16'b0000110100011010;    
    16'b0001000001001101;    
    16'b0001001001110000;    
    16'b0001001100101111;    
    16'b0001001001110000;    
    16'b0001000001001101;    
    16'b0000110100011010;    
    16'b0000100101001011;    
    16'b0000010101100111;    
    16'b0000000111101010;    
    16'b1111111100110011;    
    16'b1111110101110111;    
    16'b1111110010111100;    
    16'b1111110011011110;    
    16'b1111110110011010;    
    16'b1111111010100100;    
    16'b1111111110110000;    
    16'b0000000010000111;    
    16'b0000000100001001;    
    16'b0000000100110001;    
    16'b0000000100001101;    
    16'b0000000010111010;    
    16'b0000000001011000;    
    16'b0000000000000000;    
    16'b1111111111000011;    
    16'b1111111110100111;    
    16'b1111111110100111;    
    16'b1111111110111011;    
    16'b1111111111010110;    
    16'b1111111111110001;    
    16'b0000000000000110;    
    16'b0000000000010100;    
    16'b0000000000011010;    
    16'b0000000000011100;
    16'b0000000000000000;
    16'b0000000000000000;
    16'b0000000000000000;
    16'b0000000000000000;
  };

  always @(posedge clk) begin
    data <= rom_contents[address];
  end

endmodule
