module top_tb;

reg clk;
reg reset;
reg  signed [15:0] filter_in;
wire signed [15:0] filter_out;

reg  [11:0] filter_in_addr;
reg  filter_in_done;

reg  signed [15:0] filter_in_data_log_force [0:300]; //amostras do sinal de entrada


//  task filter_in_data_log_task; 
//  input          clk;
//  input          reset;
//  input          rdenb;   //pegar o sinal que entra no clk_enable do modulo filtro02
//  inout  [11:0]  addr;
//  output         done;
//  begin
//     if (reset == 1) 
//       addr = 0;
//     else begin
//       if (rdenb == 1) begin
//         if (addr == 300)      //testa utimo valor do verto do sinal
//           addr = addr; 
//         else
//           addr =  addr + 1; 
//       end
//     end

//     // Done Signal generation.
//     if (reset == 1)
//       done = 0; 
//     else if (addr == 300)   //testa utimo valor do verto do sinal
//       done = 1; 
//     else
//       done = 0; 
//  end
//  endtask // filter_in_data_log_task

top U1 (
	.clk (clk),
	.reset (reset),
	.filter_in (filter_in),
	.filter_out (filter_out)
);

initial
begin
	clk = 0;
	reset = 0;
	#1	reset = 1;
	#10	reset = 0;
end

always
	#5 clk = !clk;

// initial begin
// 	#10000 
// 	$fclose(f);
// 	$finish;
// end
// integer f;

// initial begin
//   f = $fopen("firpbFPGA.txt","w");
// end

// always @(posedge clk or posedge reset)
// 	filter_in_data_log_task(clk, reset, U1.SYNTHESIZED_WIRE_3, filter_in_addr, filter_in_done);

// always @ (U1.SYNTHESIZED_WIRE_3, filter_in_addr)
// begin
// 	if ( U1.SYNTHESIZED_WIRE_3 == 1) begin
//       		filter_in <= # 2 filter_in_data_log_force[filter_in_addr];
// 		$fwrite(f,"%d\n",filter_out);
//     	end
// end 

// initial //Input & Output data
//  begin
//  // Input data for filter_in_data_log
// filter_in_data_log_force[ 0   ] <=  16'b 0000000000000000 ;
// filter_in_data_log_force[ 1   ] <=  16'b 0101001111000110 ;
// filter_in_data_log_force[ 2   ] <=  16'b 0001000010111110 ;
// filter_in_data_log_force[ 3   ] <=  16'b 0001110110100011 ;
// filter_in_data_log_force[ 4   ] <=  16'b 0101100111100011 ;
// filter_in_data_log_force[ 5   ] <=  16'b 0011110110010000 ;
// filter_in_data_log_force[ 6   ] <=  16'b 0011001001000010 ;
// filter_in_data_log_force[ 7   ] <=  16'b 0001000011010011 ;
// filter_in_data_log_force[ 8   ] <= -16'b 0001111001101111 ;
// filter_in_data_log_force[ 9   ] <=  16'b 0000111011111010 ;
// filter_in_data_log_force[ 10  ] <= -16'b 0001011010100000 ;
// filter_in_data_log_force[ 11  ] <= -16'b 0111101000111110 ;
// filter_in_data_log_force[ 12  ] <= -16'b 0011011000011100 ;
// filter_in_data_log_force[ 13  ] <= -16'b 0000011001011000 ;
// filter_in_data_log_force[ 14  ] <= -16'b 0100110011011100 ;
// filter_in_data_log_force[ 15  ] <= -16'b 0010110000111110 ;
// filter_in_data_log_force[ 16  ] <=  16'b 0001001011001111 ;
// filter_in_data_log_force[ 17  ] <=  16'b 0001100010010111 ;
// filter_in_data_log_force[ 18  ] <=  16'b 0011101111001000 ;
// filter_in_data_log_force[ 19  ] <=  16'b 0010101111011001 ;
// filter_in_data_log_force[ 20  ] <=  16'b 0001111111111111 ;
// filter_in_data_log_force[ 21  ] <=  16'b 0110101111011001 ;
// filter_in_data_log_force[ 22  ] <=  16'b 0011101111001000 ;
// filter_in_data_log_force[ 23  ] <= -16'b 0010011101101000 ;
// filter_in_data_log_force[ 24  ] <=  16'b 0001001011001111 ;
// filter_in_data_log_force[ 25  ] <=  16'b 0001001111000001 ;
// filter_in_data_log_force[ 26  ] <= -16'b 0100110011011100 ;
// filter_in_data_log_force[ 27  ] <= -16'b 0100011001011000 ;
// filter_in_data_log_force[ 28  ] <= -16'b 0011011000011100 ;
// filter_in_data_log_force[ 29  ] <= -16'b 0011101000111110 ;
// filter_in_data_log_force[ 30  ] <= -16'b 0001011010100000 ;
// filter_in_data_log_force[ 31  ] <= -16'b 0011000100000101 ;
// filter_in_data_log_force[ 32  ] <= -16'b 0001111001101111 ;
// filter_in_data_log_force[ 33  ] <=  16'b 0101000011010011 ;
// filter_in_data_log_force[ 34  ] <=  16'b 0011001001000010 ;
// filter_in_data_log_force[ 35  ] <= -16'b 0000001001101111 ;
// filter_in_data_log_force[ 36  ] <=  16'b 0101100111100011 ;
// filter_in_data_log_force[ 37  ] <=  16'b 0101110110100011 ;
// filter_in_data_log_force[ 38  ] <=  16'b 0001000010111110 ;
// filter_in_data_log_force[ 39  ] <=  16'b 0001001111000110 ;
// filter_in_data_log_force[ 40  ] <=  16'b 0000000000000000 ;
// filter_in_data_log_force[ 41  ] <= -16'b 0001001111000110 ;
// filter_in_data_log_force[ 42  ] <= -16'b 0001000010111110 ;
// filter_in_data_log_force[ 43  ] <= -16'b 0101110110100011 ;
// filter_in_data_log_force[ 44  ] <= -16'b 0101100111100011 ;
// filter_in_data_log_force[ 45  ] <=  16'b 0000001001101111 ;
// filter_in_data_log_force[ 46  ] <= -16'b 0011001001000010 ;
// filter_in_data_log_force[ 47  ] <= -16'b 0101000011010011 ;
// filter_in_data_log_force[ 48  ] <=  16'b 0001111001101111 ;
// filter_in_data_log_force[ 49  ] <=  16'b 0011000100000101 ;
// filter_in_data_log_force[ 50  ] <=  16'b 0001011010100000 ;
// filter_in_data_log_force[ 51  ] <=  16'b 0011101000111110 ;
// filter_in_data_log_force[ 52  ] <=  16'b 0011011000011100 ;
// filter_in_data_log_force[ 53  ] <=  16'b 0100011001011000 ;
// filter_in_data_log_force[ 54  ] <=  16'b 0100110011011100 ;
// filter_in_data_log_force[ 55  ] <= -16'b 0001001111000001 ;
// filter_in_data_log_force[ 56  ] <= -16'b 0001001011001111 ;
// filter_in_data_log_force[ 57  ] <=  16'b 0010011101101000 ;
// filter_in_data_log_force[ 58  ] <= -16'b 0011101111001000 ;
// filter_in_data_log_force[ 59  ] <= -16'b 0110101111011001 ;
// filter_in_data_log_force[ 60  ] <= -16'b 0010000000000000 ;
// filter_in_data_log_force[ 61  ] <= -16'b 0010101111011001 ;
// filter_in_data_log_force[ 62  ] <= -16'b 0011101111001000 ;
// filter_in_data_log_force[ 63  ] <= -16'b 0001100010010111 ;
// filter_in_data_log_force[ 64  ] <= -16'b 0001001011001111 ;
// filter_in_data_log_force[ 65  ] <=  16'b 0010110000111110 ;
// filter_in_data_log_force[ 66  ] <=  16'b 0100110011011100 ;
// filter_in_data_log_force[ 67  ] <=  16'b 0000011001011000 ;
// filter_in_data_log_force[ 68  ] <=  16'b 0011011000011100 ;
// filter_in_data_log_force[ 69  ] <=  16'b 0111101000111110 ;
// filter_in_data_log_force[ 70  ] <=  16'b 0001011010100000 ;
// filter_in_data_log_force[ 71  ] <= -16'b 0000111011111010 ;
// filter_in_data_log_force[ 72  ] <=  16'b 0001111001101111 ;
// filter_in_data_log_force[ 73  ] <= -16'b 0001000011010011 ;
// filter_in_data_log_force[ 74  ] <= -16'b 0011001001000010 ;
// filter_in_data_log_force[ 75  ] <= -16'b 0011110110010000 ;
// filter_in_data_log_force[ 76  ] <= -16'b 0101100111100011 ;
// filter_in_data_log_force[ 77  ] <= -16'b 0001110110100011 ;
// filter_in_data_log_force[ 78  ] <= -16'b 0001000010111110 ;
// filter_in_data_log_force[ 79  ] <= -16'b 0101001111000110 ;
// filter_in_data_log_force[ 80  ] <=  16'b 0000000000000000 ;
// filter_in_data_log_force[ 81  ] <=  16'b 0101001111000110 ;
// filter_in_data_log_force[ 82  ] <=  16'b 0001000010111110 ;
// filter_in_data_log_force[ 83  ] <=  16'b 0001110110100011 ;
// filter_in_data_log_force[ 84  ] <=  16'b 0101100111100011 ;
// filter_in_data_log_force[ 85  ] <=  16'b 0011110110010000 ;
// filter_in_data_log_force[ 86  ] <=  16'b 0011001001000010 ;
// filter_in_data_log_force[ 87  ] <=  16'b 0001000011010011 ;
// filter_in_data_log_force[ 88  ] <= -16'b 0001111001101111 ;
// filter_in_data_log_force[ 89  ] <=  16'b 0000111011111010 ;
// filter_in_data_log_force[ 90  ] <= -16'b 0001011010100000 ;
// filter_in_data_log_force[ 91  ] <= -16'b 0111101000111110 ;
// filter_in_data_log_force[ 92  ] <= -16'b 0011011000011100 ;
// filter_in_data_log_force[ 93  ] <= -16'b 0000011001011000 ;
// filter_in_data_log_force[ 94  ] <= -16'b 0100110011011100 ;
// filter_in_data_log_force[ 95  ] <= -16'b 0010110000111110 ;
// filter_in_data_log_force[ 96  ] <=  16'b 0001001011001111 ;
// filter_in_data_log_force[ 97  ] <=  16'b 0001100010010111 ;
// filter_in_data_log_force[ 98  ] <=  16'b 0011101111001000 ;
// filter_in_data_log_force[ 99  ] <=  16'b 0010101111011001 ;
// filter_in_data_log_force[ 100 ] <=  16'b 0010000000000000 ;
// filter_in_data_log_force[ 101 ] <=  16'b 0110101111011001 ;
// filter_in_data_log_force[ 102 ] <=  16'b 0011101111001000 ;
// filter_in_data_log_force[ 103 ] <= -16'b 0010011101101000 ;
// filter_in_data_log_force[ 104 ] <=  16'b 0001001011001111 ;
// filter_in_data_log_force[ 105 ] <=  16'b 0001001111000001 ;
// filter_in_data_log_force[ 106 ] <= -16'b 0100110011011100 ;
// filter_in_data_log_force[ 107 ] <= -16'b 0100011001011000 ;
// filter_in_data_log_force[ 108 ] <= -16'b 0011011000011100 ;
// filter_in_data_log_force[ 109 ] <= -16'b 0011101000111110 ;
// filter_in_data_log_force[ 110 ] <= -16'b 0001011010100000 ;
// filter_in_data_log_force[ 111 ] <= -16'b 0011000100000101 ;
// filter_in_data_log_force[ 112 ] <= -16'b 0001111001101111 ;
// filter_in_data_log_force[ 113 ] <=  16'b 0101000011010011 ;
// filter_in_data_log_force[ 114 ] <=  16'b 0011001001000010 ;
// filter_in_data_log_force[ 115 ] <= -16'b 0000001001101111 ;
// filter_in_data_log_force[ 116 ] <=  16'b 0101100111100011 ;
// filter_in_data_log_force[ 117 ] <=  16'b 0101110110100011 ;
// filter_in_data_log_force[ 118 ] <=  16'b 0001000010111110 ;
// filter_in_data_log_force[ 119 ] <=  16'b 0001001111000110 ;
// filter_in_data_log_force[ 120 ] <=  16'b 0000000000000000 ;
// filter_in_data_log_force[ 121 ] <= -16'b 0001001111000110 ;
// filter_in_data_log_force[ 122 ] <= -16'b 0001000010111110 ;
// filter_in_data_log_force[ 123 ] <= -16'b 0101110110100011 ;
// filter_in_data_log_force[ 124 ] <= -16'b 0101100111100011 ;
// filter_in_data_log_force[ 125 ] <=  16'b 0000001001101111 ;
// filter_in_data_log_force[ 126 ] <= -16'b 0011001001000010 ;
// filter_in_data_log_force[ 127 ] <= -16'b 0101000011010011 ;
// filter_in_data_log_force[ 128 ] <=  16'b 0001111001101111 ;
// filter_in_data_log_force[ 129 ] <=  16'b 0011000100000101 ;
// filter_in_data_log_force[ 130 ] <=  16'b 0001011010100000 ;
// filter_in_data_log_force[ 131 ] <=  16'b 0011101000111110 ;
// filter_in_data_log_force[ 132 ] <=  16'b 0011011000011100 ;
// filter_in_data_log_force[ 133 ] <=  16'b 0100011001011000 ;
// filter_in_data_log_force[ 134 ] <=  16'b 0100110011011100 ;
// filter_in_data_log_force[ 135 ] <= -16'b 0001001111000001 ;
// filter_in_data_log_force[ 136 ] <= -16'b 0001001011001111 ;
// filter_in_data_log_force[ 137 ] <=  16'b 0010011101101000 ;
// filter_in_data_log_force[ 138 ] <= -16'b 0011101111001000 ;
// filter_in_data_log_force[ 139 ] <= -16'b 0110101111011001 ;
// filter_in_data_log_force[ 140 ] <= -16'b 0010000000000000 ;
// filter_in_data_log_force[ 141 ] <= -16'b 0010101111011001 ;
// filter_in_data_log_force[ 142 ] <= -16'b 0011101111001000 ;
// filter_in_data_log_force[ 143 ] <= -16'b 0001100010010111 ;
// filter_in_data_log_force[ 144 ] <= -16'b 0001001011001111 ;
// filter_in_data_log_force[ 145 ] <=  16'b 0010110000111110 ;
// filter_in_data_log_force[ 146 ] <=  16'b 0100110011011100 ;
// filter_in_data_log_force[ 147 ] <=  16'b 0000011001011000 ;
// filter_in_data_log_force[ 148 ] <=  16'b 0011011000011100 ;
// filter_in_data_log_force[ 149 ] <=  16'b 0111101000111110 ;
// filter_in_data_log_force[ 150 ] <=  16'b 0001011010100000 ;
// filter_in_data_log_force[ 151 ] <= -16'b 0000111011111010 ;
// filter_in_data_log_force[ 152 ] <=  16'b 0001111001101111 ;
// filter_in_data_log_force[ 153 ] <= -16'b 0001000011010011 ;
// filter_in_data_log_force[ 154 ] <= -16'b 0011001001000010 ;
// filter_in_data_log_force[ 155 ] <= -16'b 0011110110010000 ;
// filter_in_data_log_force[ 156 ] <= -16'b 0101100111100011 ;
// filter_in_data_log_force[ 157 ] <= -16'b 0001110110100011 ;
// filter_in_data_log_force[ 158 ] <= -16'b 0001000010111110 ;
// filter_in_data_log_force[ 159 ] <= -16'b 0101001111000110 ;
// filter_in_data_log_force[ 160 ] <=  16'b 0000000000000000 ;
// filter_in_data_log_force[ 161 ] <=  16'b 0101001111000110 ;
// filter_in_data_log_force[ 162 ] <=  16'b 0001000010111110 ;
// filter_in_data_log_force[ 163 ] <=  16'b 0001110110100011 ;
// filter_in_data_log_force[ 164 ] <=  16'b 0101100111100011 ;
// filter_in_data_log_force[ 165 ] <=  16'b 0011110110010000 ;
// filter_in_data_log_force[ 166 ] <=  16'b 0011001001000010 ;
// filter_in_data_log_force[ 167 ] <=  16'b 0001000011010011 ;
// filter_in_data_log_force[ 168 ] <= -16'b 0001111001101111 ;
// filter_in_data_log_force[ 169 ] <=  16'b 0000111011111010 ;
// filter_in_data_log_force[ 170 ] <= -16'b 0001011010100000 ;
// filter_in_data_log_force[ 171 ] <= -16'b 0111101000111110 ;
// filter_in_data_log_force[ 172 ] <= -16'b 0011011000011100 ;
// filter_in_data_log_force[ 173 ] <= -16'b 0000011001011000 ;
// filter_in_data_log_force[ 174 ] <= -16'b 0100110011011100 ;
// filter_in_data_log_force[ 175 ] <= -16'b 0010110000111110 ;
// filter_in_data_log_force[ 176 ] <=  16'b 0001001011001111 ;
// filter_in_data_log_force[ 177 ] <=  16'b 0001100010010111 ;
// filter_in_data_log_force[ 178 ] <=  16'b 0011101111001000 ;
// filter_in_data_log_force[ 179 ] <=  16'b 0010101111011001 ;
// filter_in_data_log_force[ 180 ] <=  16'b 0001111111111111 ;
// filter_in_data_log_force[ 181 ] <=  16'b 0110101111011001 ;
// filter_in_data_log_force[ 182 ] <=  16'b 0011101111001000 ;
// filter_in_data_log_force[ 183 ] <= -16'b 0010011101101000 ;
// filter_in_data_log_force[ 184 ] <=  16'b 0001001011001111 ;
// filter_in_data_log_force[ 185 ] <=  16'b 0001001111000001 ;
// filter_in_data_log_force[ 186 ] <= -16'b 0100110011011100 ;
// filter_in_data_log_force[ 187 ] <= -16'b 0100011001011000 ;
// filter_in_data_log_force[ 188 ] <= -16'b 0011011000011100 ;
// filter_in_data_log_force[ 189 ] <= -16'b 0011101000111110 ;
// filter_in_data_log_force[ 190 ] <= -16'b 0001011010100000 ;
// filter_in_data_log_force[ 191 ] <= -16'b 0011000100000101 ;
// filter_in_data_log_force[ 192 ] <= -16'b 0001111001101111 ;
// filter_in_data_log_force[ 193 ] <=  16'b 0101000011010011 ;
// filter_in_data_log_force[ 194 ] <=  16'b 0011001001000010 ;
// filter_in_data_log_force[ 195 ] <= -16'b 0000001001101111 ;
// filter_in_data_log_force[ 196 ] <=  16'b 0101100111100011 ;
// filter_in_data_log_force[ 197 ] <=  16'b 0101110110100011 ;
// filter_in_data_log_force[ 198 ] <=  16'b 0001000010111110 ;
// filter_in_data_log_force[ 199 ] <=  16'b 0001001111000110 ;
// filter_in_data_log_force[ 200 ] <=  16'b 0000000000000000 ;
// filter_in_data_log_force[ 201 ] <= -16'b 0001001111000110 ;
// filter_in_data_log_force[ 202 ] <= -16'b 0001000010111110 ;
// filter_in_data_log_force[ 203 ] <= -16'b 0101110110100011 ;
// filter_in_data_log_force[ 204 ] <= -16'b 0101100111100011 ;
// filter_in_data_log_force[ 205 ] <=  16'b 0000001001101111 ;
// filter_in_data_log_force[ 206 ] <= -16'b 0011001001000010 ;
// filter_in_data_log_force[ 207 ] <= -16'b 0101000011010011 ;
// filter_in_data_log_force[ 208 ] <=  16'b 0001111001101111 ;
// filter_in_data_log_force[ 209 ] <=  16'b 0011000100000101 ;
// filter_in_data_log_force[ 210 ] <=  16'b 0001011010100000 ;
// filter_in_data_log_force[ 211 ] <=  16'b 0011101000111110 ;
// filter_in_data_log_force[ 212 ] <=  16'b 0011011000011100 ;
// filter_in_data_log_force[ 213 ] <=  16'b 0100011001011000 ;
// filter_in_data_log_force[ 214 ] <=  16'b 0100110011011100 ;
// filter_in_data_log_force[ 215 ] <= -16'b 0001001111000001 ;
// filter_in_data_log_force[ 216 ] <= -16'b 0001001011001111 ;
// filter_in_data_log_force[ 217 ] <=  16'b 0010011101101000 ;
// filter_in_data_log_force[ 218 ] <= -16'b 0011101111001000 ;
// filter_in_data_log_force[ 219 ] <= -16'b 0110101111011001 ;
// filter_in_data_log_force[ 220 ] <= -16'b 0010000000000000 ;
// filter_in_data_log_force[ 221 ] <= -16'b 0010101111011001 ;
// filter_in_data_log_force[ 222 ] <= -16'b 0011101111001000 ;
// filter_in_data_log_force[ 223 ] <= -16'b 0001100010010111 ;
// filter_in_data_log_force[ 224 ] <= -16'b 0001001011001111 ;
// filter_in_data_log_force[ 225 ] <=  16'b 0010110000111110 ;
// filter_in_data_log_force[ 226 ] <=  16'b 0100110011011100 ;
// filter_in_data_log_force[ 227 ] <=  16'b 0000011001011000 ;
// filter_in_data_log_force[ 228 ] <=  16'b 0011011000011100 ;
// filter_in_data_log_force[ 229 ] <=  16'b 0111101000111110 ;
// filter_in_data_log_force[ 230 ] <=  16'b 0001011010100000 ;
// filter_in_data_log_force[ 231 ] <= -16'b 0000111011111010 ;
// filter_in_data_log_force[ 232 ] <=  16'b 0001111001101111 ;
// filter_in_data_log_force[ 233 ] <= -16'b 0001000011010011 ;
// filter_in_data_log_force[ 234 ] <= -16'b 0011001001000010 ;
// filter_in_data_log_force[ 235 ] <= -16'b 0011110110010000 ;
// filter_in_data_log_force[ 236 ] <= -16'b 0101100111100011 ;
// filter_in_data_log_force[ 237 ] <= -16'b 0001110110100011 ;
// filter_in_data_log_force[ 238 ] <= -16'b 0001000010111110 ;
// filter_in_data_log_force[ 239 ] <= -16'b 0101001111000110 ;
// filter_in_data_log_force[ 240 ] <=  16'b 0000000000000000 ;
// filter_in_data_log_force[ 241 ] <=  16'b 0101001111000110 ;
// filter_in_data_log_force[ 242 ] <=  16'b 0001000010111110 ;
// filter_in_data_log_force[ 243 ] <=  16'b 0001110110100011 ;
// filter_in_data_log_force[ 244 ] <=  16'b 0101100111100011 ;
// filter_in_data_log_force[ 245 ] <=  16'b 0011110110010000 ;
// filter_in_data_log_force[ 246 ] <=  16'b 0011001001000010 ;
// filter_in_data_log_force[ 247 ] <=  16'b 0001000011010011 ;
// filter_in_data_log_force[ 248 ] <= -16'b 0001111001101111 ;
// filter_in_data_log_force[ 249 ] <=  16'b 0000111011111010 ;
// filter_in_data_log_force[ 250 ] <= -16'b 0001011010100000 ;
// filter_in_data_log_force[ 251 ] <= -16'b 0111101000111110 ;
// filter_in_data_log_force[ 252 ] <= -16'b 0011011000011100 ;
// filter_in_data_log_force[ 253 ] <= -16'b 0000011001011000 ;
// filter_in_data_log_force[ 254 ] <= -16'b 0100110011011100 ;
// filter_in_data_log_force[ 255 ] <= -16'b 0010110000111110 ;
// filter_in_data_log_force[ 256 ] <=  16'b 0001001011001111 ;
// filter_in_data_log_force[ 257 ] <=  16'b 0001100010010111 ;
// filter_in_data_log_force[ 258 ] <=  16'b 0011101111001000 ;
// filter_in_data_log_force[ 259 ] <=  16'b 0010101111011001 ;
// filter_in_data_log_force[ 260 ] <=  16'b 0001111111111111 ;
// filter_in_data_log_force[ 261 ] <=  16'b 0110101111011001 ;
// filter_in_data_log_force[ 262 ] <=  16'b 0011101111001000 ;
// filter_in_data_log_force[ 263 ] <= -16'b 0010011101101000 ;
// filter_in_data_log_force[ 264 ] <=  16'b 0001001011001111 ;
// filter_in_data_log_force[ 265 ] <=  16'b 0001001111000001 ;
// filter_in_data_log_force[ 266 ] <= -16'b 0100110011011100 ;
// filter_in_data_log_force[ 267 ] <= -16'b 0100011001011000 ;
// filter_in_data_log_force[ 268 ] <= -16'b 0011011000011100 ;
// filter_in_data_log_force[ 269 ] <= -16'b 0011101000111110 ;
// filter_in_data_log_force[ 270 ] <= -16'b 0001011010100000 ;
// filter_in_data_log_force[ 271 ] <= -16'b 0011000100000101 ;
// filter_in_data_log_force[ 272 ] <= -16'b 0001111001101111 ;
// filter_in_data_log_force[ 273 ] <=  16'b 0101000011010011 ;
// filter_in_data_log_force[ 274 ] <=  16'b 0011001001000010 ;
// filter_in_data_log_force[ 275 ] <= -16'b 0000001001101111 ;
// filter_in_data_log_force[ 276 ] <=  16'b 0101100111100011 ;
// filter_in_data_log_force[ 277 ] <=  16'b 0101110110100011 ;
// filter_in_data_log_force[ 278 ] <=  16'b 0001000010111110 ;
// filter_in_data_log_force[ 279 ] <=  16'b 0001001111000110 ;
// filter_in_data_log_force[ 280 ] <=  16'b 0000000000000000 ;
// filter_in_data_log_force[ 281 ] <= -16'b 0001001111000110 ;
// filter_in_data_log_force[ 282 ] <= -16'b 0001000010111110 ;
// filter_in_data_log_force[ 283 ] <= -16'b 0101110110100011 ;
// filter_in_data_log_force[ 284 ] <= -16'b 0101100111100011 ;
// filter_in_data_log_force[ 285 ] <=  16'b 0000001001101111 ;
// filter_in_data_log_force[ 286 ] <= -16'b 0011001001000010 ;
// filter_in_data_log_force[ 287 ] <= -16'b 0101000011010011 ;
// filter_in_data_log_force[ 288 ] <=  16'b 0001111001101111 ;
// filter_in_data_log_force[ 289 ] <=  16'b 0011000100000101 ;
// filter_in_data_log_force[ 290 ] <=  16'b 0001011010100000 ;
// filter_in_data_log_force[ 291 ] <=  16'b 0011101000111110 ;
// filter_in_data_log_force[ 292 ] <=  16'b 0011011000011100 ;
// filter_in_data_log_force[ 293 ] <=  16'b 0100011001011000 ;
// filter_in_data_log_force[ 294 ] <=  16'b 0100110011011100 ;
// filter_in_data_log_force[ 295 ] <= -16'b 0001001111000001 ;
// filter_in_data_log_force[ 296 ] <= -16'b 0001001011001111 ;
// filter_in_data_log_force[ 297 ] <=  16'b 0010011101101000 ;
// filter_in_data_log_force[ 298 ] <= -16'b 0011101111001000 ;
// filter_in_data_log_force[ 299 ] <= -16'b 0110101111011001 ;
// end 
endmodule 
